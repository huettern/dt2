library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
	port (
		rst_n : in std_ulogic;
		btn_n : in std_ulogic;
		clk : in std_ulogic;
		hex_n : out std_ulogic_vector
	);
end entity top;

architecture structural of top is

begin

end architecture structural;
